
`define A
`define B
`define C
`ifdef X
1
2
`endif
4

6

