
`define A
`define B
`define C

1
2
4

6

